module SON3 (
    input  wire                clk            ,
	input  wire                rst_n          ,
	input  wire  [3:0]         cfg_of_son3    ,
	input  wire  [15:0]        dout_of_son1_1 ,
	input  wire  [15:0]        dout_of_son1_2 ,
	input  wire  [15:0]        dout_of_son2 ,
	output wire  [15:0]        dout_of_son3


);

endmodule
